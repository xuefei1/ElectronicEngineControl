// niosII_system.v

// Generated using ACDS version 12.1sp1 243 at 2017.03.17.16:47:28

`timescale 1 ps / 1 ps
module niosII_system (
		output wire        altpll_0_c0_out,                         //                       altpll_0_c0.clk
		input  wire        rs232_0_external_interface_RXD,          //        rs232_0_external_interface.RXD
		output wire        rs232_0_external_interface_TXD,          //                                  .TXD
		output wire        pwm_generator_0_pwm_out_export,          //           pwm_generator_0_pwm_out.export
		output wire        phasedone_from_the_altpll_0,             //        altpll_0_phasedone_conduit.export
		input  wire        reset_n,                                 //                clk_0_clk_in_reset.reset_n
		input  wire        in_port_to_the_switch,                   //        switch_external_connection.export
		output wire [12:0] sdram_0_wire_addr,                       //                      sdram_0_wire.addr
		output wire [1:0]  sdram_0_wire_ba,                         //                                  .ba
		output wire        sdram_0_wire_cas_n,                      //                                  .cas_n
		output wire        sdram_0_wire_cke,                        //                                  .cke
		output wire        sdram_0_wire_cs_n,                       //                                  .cs_n
		inout  wire [15:0] sdram_0_wire_dq,                         //                                  .dq
		output wire [1:0]  sdram_0_wire_dqm,                        //                                  .dqm
		output wire        sdram_0_wire_ras_n,                      //                                  .ras_n
		output wire        sdram_0_wire_we_n,                       //                                  .we_n
		output wire [7:0]  out_port_from_the_green_leds,            //    green_leds_external_connection.export
		output wire [7:0]  solenoid_out_external_connection_export, //  solenoid_out_external_connection.export
		input  wire        areset_to_the_altpll_0,                  //           altpll_0_areset_conduit.export
		output wire        locked_from_the_altpll_0,                //           altpll_0_locked_conduit.export
		input  wire        clk_0,                                   //                      clk_0_clk_in.clk
		output wire        adc_sclk_from_the_de0_nano_adc_0,        // de0_nano_adc_0_external_interface.sclk
		output wire        adc_cs_n_from_the_de0_nano_adc_0,        //                                  .cs_n
		input  wire        adc_dout_to_the_de0_nano_adc_0,          //                                  .dout
		output wire        adc_din_from_the_de0_nano_adc_0,         //                                  .din
		input  wire [7:0]  buttons_external_connection_export       //       buttons_external_connection.export
	);

	wire          altpll_0_c1_clk;                                                                                           // altpll_0:c1 -> [addr_router:clk, addr_router_001:clk, burst_adapter:clk, burst_adapter_001:clk, buttons:clk, buttons_s1_translator:clk, buttons_s1_translator_avalon_universal_slave_0_agent:clk, buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, crosser:in_clk, crosser_001:out_clk, de0_nano_adc_0:clock, de0_nano_adc_0_adc_slave_translator:clk, de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:clk, de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, green_leds:clk, green_leds_s1_translator:clk, green_leds_s1_translator_avalon_universal_slave_0_agent:clk, green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, irq_mapper:clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, nios2_0:clk, nios2_0_data_master_translator:clk, nios2_0_data_master_translator_avalon_universal_master_0_agent:clk, nios2_0_instruction_master_translator:clk, nios2_0_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_0_jtag_debug_module_translator:clk, nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2_0:clk, onchip_memory2_0_s1_translator:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pwm_generator_0:clock, pwm_generator_0_avalon_slave_control_translator:clk, pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:clk, pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pwm_generator_0_avalon_slave_duty_translator:clk, pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:clk, pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pwm_generator_0_avalon_slave_period_translator:clk, pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:clk, pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rs232_0:clk, rs232_0_avalon_rs232_slave_translator:clk, rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:clk, rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, sdram_0:clk, sdram_0_s1_translator:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, solenoid_out:clk, solenoid_out_s1_translator:clk, solenoid_out_s1_translator_avalon_universal_slave_0_agent:clk, solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, switch:clk, switch_s1_translator:clk, switch_s1_translator_avalon_universal_slave_0_agent:clk, switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sys_clk_timer:clk, sys_clk_timer_s1_translator:clk, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:clk, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sysid_qsys_0:clock, sysid_qsys_0_control_slave_translator:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timestamp_timer:clk, timestamp_timer_s1_translator:clk, timestamp_timer_s1_translator_avalon_universal_slave_0_agent:clk, timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk]
	wire          nios2_0_jtag_debug_module_reset_reset;                                                                     // nios2_0:jtag_debug_module_resetrequest -> [burst_adapter:reset, burst_adapter_001:reset, buttons:reset_n, buttons_s1_translator:reset, buttons_s1_translator_avalon_universal_slave_0_agent:reset, buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_mux_002:reset, id_router_002:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, pwm_generator_0:reset, pwm_generator_0_avalon_slave_control_translator:reset, pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:reset, pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pwm_generator_0_avalon_slave_duty_translator:reset, pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:reset, pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pwm_generator_0_avalon_slave_period_translator:reset, pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:reset, pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rs232_0:reset, rs232_0_avalon_rs232_slave_translator:reset, rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:reset, rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rst_controller:reset_in1, rst_controller_001:reset_in1, sdram_0:reset_n, sdram_0_s1_translator:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, solenoid_out:reset_n, solenoid_out_s1_translator:reset, solenoid_out_s1_translator_avalon_universal_slave_0_agent:reset, solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timestamp_timer:reset_n, timestamp_timer_s1_translator:reset, timestamp_timer_s1_translator_avalon_universal_slave_0_agent:reset, timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          nios2_0_instruction_master_waitrequest;                                                                    // nios2_0_instruction_master_translator:av_waitrequest -> nios2_0:i_waitrequest
	wire   [26:0] nios2_0_instruction_master_address;                                                                        // nios2_0:i_address -> nios2_0_instruction_master_translator:av_address
	wire          nios2_0_instruction_master_read;                                                                           // nios2_0:i_read -> nios2_0_instruction_master_translator:av_read
	wire   [31:0] nios2_0_instruction_master_readdata;                                                                       // nios2_0_instruction_master_translator:av_readdata -> nios2_0:i_readdata
	wire          nios2_0_data_master_waitrequest;                                                                           // nios2_0_data_master_translator:av_waitrequest -> nios2_0:d_waitrequest
	wire   [31:0] nios2_0_data_master_writedata;                                                                             // nios2_0:d_writedata -> nios2_0_data_master_translator:av_writedata
	wire   [26:0] nios2_0_data_master_address;                                                                               // nios2_0:d_address -> nios2_0_data_master_translator:av_address
	wire          nios2_0_data_master_write;                                                                                 // nios2_0:d_write -> nios2_0_data_master_translator:av_write
	wire          nios2_0_data_master_read;                                                                                  // nios2_0:d_read -> nios2_0_data_master_translator:av_read
	wire   [31:0] nios2_0_data_master_readdata;                                                                              // nios2_0_data_master_translator:av_readdata -> nios2_0:d_readdata
	wire          nios2_0_data_master_debugaccess;                                                                           // nios2_0:jtag_debug_module_debugaccess_to_roms -> nios2_0_data_master_translator:av_debugaccess
	wire    [3:0] nios2_0_data_master_byteenable;                                                                            // nios2_0:d_byteenable -> nios2_0_data_master_translator:av_byteenable
	wire   [31:0] nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                        // nios2_0_jtag_debug_module_translator:av_writedata -> nios2_0:jtag_debug_module_writedata
	wire    [8:0] nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                          // nios2_0_jtag_debug_module_translator:av_address -> nios2_0:jtag_debug_module_address
	wire          nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                                       // nios2_0_jtag_debug_module_translator:av_chipselect -> nios2_0:jtag_debug_module_select
	wire          nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                            // nios2_0_jtag_debug_module_translator:av_write -> nios2_0:jtag_debug_module_write
	wire   [31:0] nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                         // nios2_0:jtag_debug_module_readdata -> nios2_0_jtag_debug_module_translator:av_readdata
	wire          nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                                    // nios2_0_jtag_debug_module_translator:av_begintransfer -> nios2_0:jtag_debug_module_begintransfer
	wire          nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                      // nios2_0_jtag_debug_module_translator:av_debugaccess -> nios2_0:jtag_debug_module_debugaccess
	wire    [3:0] nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                       // nios2_0_jtag_debug_module_translator:av_byteenable -> nios2_0:jtag_debug_module_byteenable
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                              // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire   [11:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                                // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                             // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                                  // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                                  // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                               // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                             // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire          sdram_0_s1_translator_avalon_anti_slave_0_waitrequest;                                                     // sdram_0:za_waitrequest -> sdram_0_s1_translator:av_waitrequest
	wire   [15:0] sdram_0_s1_translator_avalon_anti_slave_0_writedata;                                                       // sdram_0_s1_translator:av_writedata -> sdram_0:az_data
	wire   [23:0] sdram_0_s1_translator_avalon_anti_slave_0_address;                                                         // sdram_0_s1_translator:av_address -> sdram_0:az_addr
	wire          sdram_0_s1_translator_avalon_anti_slave_0_chipselect;                                                      // sdram_0_s1_translator:av_chipselect -> sdram_0:az_cs
	wire          sdram_0_s1_translator_avalon_anti_slave_0_write;                                                           // sdram_0_s1_translator:av_write -> sdram_0:az_wr_n
	wire          sdram_0_s1_translator_avalon_anti_slave_0_read;                                                            // sdram_0_s1_translator:av_read -> sdram_0:az_rd_n
	wire   [15:0] sdram_0_s1_translator_avalon_anti_slave_0_readdata;                                                        // sdram_0:za_data -> sdram_0_s1_translator:av_readdata
	wire          sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid;                                                   // sdram_0:za_valid -> sdram_0_s1_translator:av_readdatavalid
	wire    [1:0] sdram_0_s1_translator_avalon_anti_slave_0_byteenable;                                                      // sdram_0_s1_translator:av_byteenable -> sdram_0:az_be_n
	wire    [0:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address;                                         // sysid_qsys_0_control_slave_translator:av_address -> sysid_qsys_0:address
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata;                                        // sysid_qsys_0:readdata -> sysid_qsys_0_control_slave_translator:av_readdata
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata;                                                 // sys_clk_timer_s1_translator:av_writedata -> sys_clk_timer:writedata
	wire    [2:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_address;                                                   // sys_clk_timer_s1_translator:av_address -> sys_clk_timer:address
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect;                                                // sys_clk_timer_s1_translator:av_chipselect -> sys_clk_timer:chipselect
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_write;                                                     // sys_clk_timer_s1_translator:av_write -> sys_clk_timer:write_n
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata;                                                  // sys_clk_timer:readdata -> sys_clk_timer_s1_translator:av_readdata
	wire   [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata;                                               // altpll_0_pll_slave_translator:av_writedata -> altpll_0:writedata
	wire    [1:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_address;                                                 // altpll_0_pll_slave_translator:av_address -> altpll_0:address
	wire          altpll_0_pll_slave_translator_avalon_anti_slave_0_write;                                                   // altpll_0_pll_slave_translator:av_write -> altpll_0:write
	wire          altpll_0_pll_slave_translator_avalon_anti_slave_0_read;                                                    // altpll_0_pll_slave_translator:av_read -> altpll_0:read
	wire   [31:0] altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata;                                                // altpll_0:readdata -> altpll_0_pll_slave_translator:av_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                  // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                    // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire    [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                      // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                        // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                         // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                     // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] green_leds_s1_translator_avalon_anti_slave_0_writedata;                                                    // green_leds_s1_translator:av_writedata -> green_leds:writedata
	wire    [1:0] green_leds_s1_translator_avalon_anti_slave_0_address;                                                      // green_leds_s1_translator:av_address -> green_leds:address
	wire          green_leds_s1_translator_avalon_anti_slave_0_chipselect;                                                   // green_leds_s1_translator:av_chipselect -> green_leds:chipselect
	wire          green_leds_s1_translator_avalon_anti_slave_0_write;                                                        // green_leds_s1_translator:av_write -> green_leds:write_n
	wire   [31:0] green_leds_s1_translator_avalon_anti_slave_0_readdata;                                                     // green_leds:readdata -> green_leds_s1_translator:av_readdata
	wire    [1:0] switch_s1_translator_avalon_anti_slave_0_address;                                                          // switch_s1_translator:av_address -> switch:address
	wire   [31:0] switch_s1_translator_avalon_anti_slave_0_readdata;                                                         // switch:readdata -> switch_s1_translator:av_readdata
	wire          de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_waitrequest;                                       // de0_nano_adc_0:waitrequest -> de0_nano_adc_0_adc_slave_translator:av_waitrequest
	wire   [31:0] de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_writedata;                                         // de0_nano_adc_0_adc_slave_translator:av_writedata -> de0_nano_adc_0:writedata
	wire    [2:0] de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_address;                                           // de0_nano_adc_0_adc_slave_translator:av_address -> de0_nano_adc_0:address
	wire          de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_write;                                             // de0_nano_adc_0_adc_slave_translator:av_write -> de0_nano_adc_0:write
	wire          de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_read;                                              // de0_nano_adc_0_adc_slave_translator:av_read -> de0_nano_adc_0:read
	wire   [31:0] de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_readdata;                                          // de0_nano_adc_0:readdata -> de0_nano_adc_0_adc_slave_translator:av_readdata
	wire   [31:0] rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata;                                       // rs232_0_avalon_rs232_slave_translator:av_writedata -> rs232_0:writedata
	wire    [0:0] rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_address;                                         // rs232_0_avalon_rs232_slave_translator:av_address -> rs232_0:address
	wire          rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect;                                      // rs232_0_avalon_rs232_slave_translator:av_chipselect -> rs232_0:chipselect
	wire          rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_write;                                           // rs232_0_avalon_rs232_slave_translator:av_write -> rs232_0:write
	wire          rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_read;                                            // rs232_0_avalon_rs232_slave_translator:av_read -> rs232_0:read
	wire   [31:0] rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata;                                        // rs232_0:readdata -> rs232_0_avalon_rs232_slave_translator:av_readdata
	wire    [3:0] rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable;                                      // rs232_0_avalon_rs232_slave_translator:av_byteenable -> rs232_0:byteenable
	wire   [15:0] timestamp_timer_s1_translator_avalon_anti_slave_0_writedata;                                               // timestamp_timer_s1_translator:av_writedata -> timestamp_timer:writedata
	wire    [2:0] timestamp_timer_s1_translator_avalon_anti_slave_0_address;                                                 // timestamp_timer_s1_translator:av_address -> timestamp_timer:address
	wire          timestamp_timer_s1_translator_avalon_anti_slave_0_chipselect;                                              // timestamp_timer_s1_translator:av_chipselect -> timestamp_timer:chipselect
	wire          timestamp_timer_s1_translator_avalon_anti_slave_0_write;                                                   // timestamp_timer_s1_translator:av_write -> timestamp_timer:write_n
	wire   [15:0] timestamp_timer_s1_translator_avalon_anti_slave_0_readdata;                                                // timestamp_timer:readdata -> timestamp_timer_s1_translator:av_readdata
	wire   [31:0] pwm_generator_0_avalon_slave_period_translator_avalon_anti_slave_0_writedata;                              // pwm_generator_0_avalon_slave_period_translator:av_writedata -> pwm_generator_0:period_in
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_anti_slave_0_write;                                  // pwm_generator_0_avalon_slave_period_translator:av_write -> pwm_generator_0:write_en_period
	wire   [31:0] pwm_generator_0_avalon_slave_duty_translator_avalon_anti_slave_0_writedata;                                // pwm_generator_0_avalon_slave_duty_translator:av_writedata -> pwm_generator_0:duty_in
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_anti_slave_0_write;                                    // pwm_generator_0_avalon_slave_duty_translator:av_write -> pwm_generator_0:write_en_duty
	wire   [31:0] buttons_s1_translator_avalon_anti_slave_0_writedata;                                                       // buttons_s1_translator:av_writedata -> buttons:writedata
	wire    [1:0] buttons_s1_translator_avalon_anti_slave_0_address;                                                         // buttons_s1_translator:av_address -> buttons:address
	wire          buttons_s1_translator_avalon_anti_slave_0_chipselect;                                                      // buttons_s1_translator:av_chipselect -> buttons:chipselect
	wire          buttons_s1_translator_avalon_anti_slave_0_write;                                                           // buttons_s1_translator:av_write -> buttons:write_n
	wire   [31:0] buttons_s1_translator_avalon_anti_slave_0_readdata;                                                        // buttons:readdata -> buttons_s1_translator:av_readdata
	wire   [31:0] solenoid_out_s1_translator_avalon_anti_slave_0_writedata;                                                  // solenoid_out_s1_translator:av_writedata -> solenoid_out:writedata
	wire    [2:0] solenoid_out_s1_translator_avalon_anti_slave_0_address;                                                    // solenoid_out_s1_translator:av_address -> solenoid_out:address
	wire          solenoid_out_s1_translator_avalon_anti_slave_0_chipselect;                                                 // solenoid_out_s1_translator:av_chipselect -> solenoid_out:chipselect
	wire          solenoid_out_s1_translator_avalon_anti_slave_0_write;                                                      // solenoid_out_s1_translator:av_write -> solenoid_out:write_n
	wire   [31:0] solenoid_out_s1_translator_avalon_anti_slave_0_readdata;                                                   // solenoid_out:readdata -> solenoid_out_s1_translator:av_readdata
	wire    [7:0] pwm_generator_0_avalon_slave_control_translator_avalon_anti_slave_0_writedata;                             // pwm_generator_0_avalon_slave_control_translator:av_writedata -> pwm_generator_0:control_in
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_anti_slave_0_write;                                 // pwm_generator_0_avalon_slave_control_translator:av_write -> pwm_generator_0:write_en_control
	wire          nios2_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                               // nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_0_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_0_instruction_master_translator_avalon_universal_master_0_burstcount;                                // nios2_0_instruction_master_translator:uav_burstcount -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_0_instruction_master_translator_avalon_universal_master_0_writedata;                                 // nios2_0_instruction_master_translator:uav_writedata -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [26:0] nios2_0_instruction_master_translator_avalon_universal_master_0_address;                                   // nios2_0_instruction_master_translator:uav_address -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_0_instruction_master_translator_avalon_universal_master_0_lock;                                      // nios2_0_instruction_master_translator:uav_lock -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_0_instruction_master_translator_avalon_universal_master_0_write;                                     // nios2_0_instruction_master_translator:uav_write -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_0_instruction_master_translator_avalon_universal_master_0_read;                                      // nios2_0_instruction_master_translator:uav_read -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_0_instruction_master_translator_avalon_universal_master_0_readdata;                                  // nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_0_instruction_master_translator:uav_readdata
	wire          nios2_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                               // nios2_0_instruction_master_translator:uav_debugaccess -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_0_instruction_master_translator_avalon_universal_master_0_byteenable;                                // nios2_0_instruction_master_translator:uav_byteenable -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                             // nios2_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_0_instruction_master_translator:uav_readdatavalid
	wire          nios2_0_data_master_translator_avalon_universal_master_0_waitrequest;                                      // nios2_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_0_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_0_data_master_translator_avalon_universal_master_0_burstcount;                                       // nios2_0_data_master_translator:uav_burstcount -> nios2_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_0_data_master_translator_avalon_universal_master_0_writedata;                                        // nios2_0_data_master_translator:uav_writedata -> nios2_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [26:0] nios2_0_data_master_translator_avalon_universal_master_0_address;                                          // nios2_0_data_master_translator:uav_address -> nios2_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_0_data_master_translator_avalon_universal_master_0_lock;                                             // nios2_0_data_master_translator:uav_lock -> nios2_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_0_data_master_translator_avalon_universal_master_0_write;                                            // nios2_0_data_master_translator:uav_write -> nios2_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_0_data_master_translator_avalon_universal_master_0_read;                                             // nios2_0_data_master_translator:uav_read -> nios2_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_0_data_master_translator_avalon_universal_master_0_readdata;                                         // nios2_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_0_data_master_translator:uav_readdata
	wire          nios2_0_data_master_translator_avalon_universal_master_0_debugaccess;                                      // nios2_0_data_master_translator:uav_debugaccess -> nios2_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_0_data_master_translator_avalon_universal_master_0_byteenable;                                       // nios2_0_data_master_translator:uav_byteenable -> nios2_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_0_data_master_translator_avalon_universal_master_0_readdatavalid;                                    // nios2_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_0_data_master_translator:uav_readdatavalid
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // nios2_0_jtag_debug_module_translator:uav_waitrequest -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_0_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                          // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_0_jtag_debug_module_translator:uav_writedata
	wire   [26:0] nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                            // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_0_jtag_debug_module_translator:uav_address
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                              // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_0_jtag_debug_module_translator:uav_write
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                               // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_0_jtag_debug_module_translator:uav_lock
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                               // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_0_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                           // nios2_0_jtag_debug_module_translator:uav_readdata -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // nios2_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_0_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_0_jtag_debug_module_translator:uav_byteenable
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                        // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire   [26:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // sdram_0_s1_translator:uav_waitrequest -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_s1_translator:uav_burstcount
	wire   [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_s1_translator:uav_writedata
	wire   [26:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_s1_translator:uav_address
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_s1_translator:uav_write
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_s1_translator:uav_lock
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_s1_translator:uav_read
	wire   [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // sdram_0_s1_translator:uav_readdata -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // sdram_0_s1_translator:uav_readdatavalid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_s1_translator:uav_debugaccess
	wire    [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_s1_translator:uav_byteenable
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [86:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [86:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // sysid_qsys_0_control_slave_translator:uav_waitrequest -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_0_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_0_control_slave_translator:uav_writedata
	wire   [26:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_0_control_slave_translator:uav_address
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_0_control_slave_translator:uav_write
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_0_control_slave_translator:uav_lock
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_0_control_slave_translator:uav_read
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // sysid_qsys_0_control_slave_translator:uav_readdata -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // sysid_qsys_0_control_slave_translator:uav_readdatavalid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_0_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_0_control_slave_translator:uav_byteenable
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // sys_clk_timer_s1_translator:uav_waitrequest -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sys_clk_timer_s1_translator:uav_burstcount
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sys_clk_timer_s1_translator:uav_writedata
	wire   [26:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sys_clk_timer_s1_translator:uav_address
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sys_clk_timer_s1_translator:uav_write
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sys_clk_timer_s1_translator:uav_lock
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sys_clk_timer_s1_translator:uav_read
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // sys_clk_timer_s1_translator:uav_readdata -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // sys_clk_timer_s1_translator:uav_readdatavalid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sys_clk_timer_s1_translator:uav_debugaccess
	wire    [3:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sys_clk_timer_s1_translator:uav_byteenable
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // altpll_0_pll_slave_translator:uav_waitrequest -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> altpll_0_pll_slave_translator:uav_burstcount
	wire   [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> altpll_0_pll_slave_translator:uav_writedata
	wire   [26:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> altpll_0_pll_slave_translator:uav_address
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                                     // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> altpll_0_pll_slave_translator:uav_write
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> altpll_0_pll_slave_translator:uav_lock
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> altpll_0_pll_slave_translator:uav_read
	wire   [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // altpll_0_pll_slave_translator:uav_readdata -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // altpll_0_pll_slave_translator:uav_readdatavalid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> altpll_0_pll_slave_translator:uav_debugaccess
	wire    [3:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> altpll_0_pll_slave_translator:uav_byteenable
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                               // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                          // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire   [26:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                       // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // green_leds_s1_translator:uav_waitrequest -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> green_leds_s1_translator:uav_burstcount
	wire   [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> green_leds_s1_translator:uav_writedata
	wire   [26:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_address -> green_leds_s1_translator:uav_address
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_write -> green_leds_s1_translator:uav_write
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_lock -> green_leds_s1_translator:uav_lock
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_read -> green_leds_s1_translator:uav_read
	wire   [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // green_leds_s1_translator:uav_readdata -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // green_leds_s1_translator:uav_readdatavalid -> green_leds_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> green_leds_s1_translator:uav_debugaccess
	wire    [3:0] green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // green_leds_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> green_leds_s1_translator:uav_byteenable
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // green_leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // switch_s1_translator:uav_waitrequest -> switch_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // switch_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch_s1_translator:uav_burstcount
	wire   [31:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // switch_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch_s1_translator:uav_writedata
	wire   [26:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_address;                                            // switch_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch_s1_translator:uav_address
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_write;                                              // switch_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch_s1_translator:uav_write
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                               // switch_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch_s1_translator:uav_lock
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_read;                                               // switch_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch_s1_translator:uav_read
	wire   [31:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // switch_s1_translator:uav_readdata -> switch_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // switch_s1_translator:uav_readdatavalid -> switch_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // switch_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch_s1_translator:uav_debugaccess
	wire    [3:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // switch_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch_s1_translator:uav_byteenable
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // de0_nano_adc_0_adc_slave_translator:uav_waitrequest -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> de0_nano_adc_0_adc_slave_translator:uav_burstcount
	wire   [31:0] de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                           // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> de0_nano_adc_0_adc_slave_translator:uav_writedata
	wire   [26:0] de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_address;                             // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_address -> de0_nano_adc_0_adc_slave_translator:uav_address
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_write;                               // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_write -> de0_nano_adc_0_adc_slave_translator:uav_write
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_lock -> de0_nano_adc_0_adc_slave_translator:uav_lock
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_read;                                // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_read -> de0_nano_adc_0_adc_slave_translator:uav_read
	wire   [31:0] de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                            // de0_nano_adc_0_adc_slave_translator:uav_readdata -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // de0_nano_adc_0_adc_slave_translator:uav_readdatavalid -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> de0_nano_adc_0_adc_slave_translator:uav_debugaccess
	wire    [3:0] de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> de0_nano_adc_0_adc_slave_translator:uav_byteenable
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                         // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // rs232_0_avalon_rs232_slave_translator:uav_waitrequest -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> rs232_0_avalon_rs232_slave_translator:uav_burstcount
	wire   [31:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                         // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> rs232_0_avalon_rs232_slave_translator:uav_writedata
	wire   [26:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address;                           // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_address -> rs232_0_avalon_rs232_slave_translator:uav_address
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write;                             // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_write -> rs232_0_avalon_rs232_slave_translator:uav_write
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock;                              // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_lock -> rs232_0_avalon_rs232_slave_translator:uav_lock
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read;                              // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_read -> rs232_0_avalon_rs232_slave_translator:uav_read
	wire   [31:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                          // rs232_0_avalon_rs232_slave_translator:uav_readdata -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // rs232_0_avalon_rs232_slave_translator:uav_readdatavalid -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> rs232_0_avalon_rs232_slave_translator:uav_debugaccess
	wire    [3:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> rs232_0_avalon_rs232_slave_translator:uav_byteenable
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                       // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // timestamp_timer_s1_translator:uav_waitrequest -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timestamp_timer_s1_translator:uav_burstcount
	wire   [31:0] timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timestamp_timer_s1_translator:uav_writedata
	wire   [26:0] timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> timestamp_timer_s1_translator:uav_address
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> timestamp_timer_s1_translator:uav_write
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timestamp_timer_s1_translator:uav_lock
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> timestamp_timer_s1_translator:uav_read
	wire   [31:0] timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // timestamp_timer_s1_translator:uav_readdata -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // timestamp_timer_s1_translator:uav_readdatavalid -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timestamp_timer_s1_translator:uav_debugaccess
	wire    [3:0] timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timestamp_timer_s1_translator:uav_byteenable
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // pwm_generator_0_avalon_slave_period_translator:uav_waitrequest -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_burstcount;               // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_burstcount -> pwm_generator_0_avalon_slave_period_translator:uav_burstcount
	wire   [31:0] pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_writedata;                // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_writedata -> pwm_generator_0_avalon_slave_period_translator:uav_writedata
	wire   [26:0] pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_address;                  // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_address -> pwm_generator_0_avalon_slave_period_translator:uav_address
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_write;                    // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_write -> pwm_generator_0_avalon_slave_period_translator:uav_write
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_lock;                     // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_lock -> pwm_generator_0_avalon_slave_period_translator:uav_lock
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_read;                     // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_read -> pwm_generator_0_avalon_slave_period_translator:uav_read
	wire   [31:0] pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_readdata;                 // pwm_generator_0_avalon_slave_period_translator:uav_readdata -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // pwm_generator_0_avalon_slave_period_translator:uav_readdatavalid -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pwm_generator_0_avalon_slave_period_translator:uav_debugaccess
	wire    [3:0] pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_byteenable;               // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:m0_byteenable -> pwm_generator_0_avalon_slave_period_translator:uav_byteenable
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_valid;             // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rf_source_valid -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_data;              // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rf_source_data -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_ready;             // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // pwm_generator_0_avalon_slave_duty_translator:uav_waitrequest -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_burstcount -> pwm_generator_0_avalon_slave_duty_translator:uav_burstcount
	wire   [31:0] pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_writedata;                  // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_writedata -> pwm_generator_0_avalon_slave_duty_translator:uav_writedata
	wire   [26:0] pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_address;                    // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_address -> pwm_generator_0_avalon_slave_duty_translator:uav_address
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_write;                      // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_write -> pwm_generator_0_avalon_slave_duty_translator:uav_write
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_lock;                       // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_lock -> pwm_generator_0_avalon_slave_duty_translator:uav_lock
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_read;                       // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_read -> pwm_generator_0_avalon_slave_duty_translator:uav_read
	wire   [31:0] pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_readdata;                   // pwm_generator_0_avalon_slave_duty_translator:uav_readdata -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // pwm_generator_0_avalon_slave_duty_translator:uav_readdatavalid -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pwm_generator_0_avalon_slave_duty_translator:uav_debugaccess
	wire    [3:0] pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:m0_byteenable -> pwm_generator_0_avalon_slave_duty_translator:uav_byteenable
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_valid;               // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rf_source_valid -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_data;                // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rf_source_data -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_ready;               // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // buttons_s1_translator:uav_waitrequest -> buttons_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] buttons_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // buttons_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> buttons_s1_translator:uav_burstcount
	wire   [31:0] buttons_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // buttons_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> buttons_s1_translator:uav_writedata
	wire   [26:0] buttons_s1_translator_avalon_universal_slave_0_agent_m0_address;                                           // buttons_s1_translator_avalon_universal_slave_0_agent:m0_address -> buttons_s1_translator:uav_address
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_m0_write;                                             // buttons_s1_translator_avalon_universal_slave_0_agent:m0_write -> buttons_s1_translator:uav_write
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                              // buttons_s1_translator_avalon_universal_slave_0_agent:m0_lock -> buttons_s1_translator:uav_lock
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_m0_read;                                              // buttons_s1_translator_avalon_universal_slave_0_agent:m0_read -> buttons_s1_translator:uav_read
	wire   [31:0] buttons_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // buttons_s1_translator:uav_readdata -> buttons_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // buttons_s1_translator:uav_readdatavalid -> buttons_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // buttons_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> buttons_s1_translator:uav_debugaccess
	wire    [3:0] buttons_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // buttons_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> buttons_s1_translator:uav_byteenable
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // buttons_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // buttons_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // buttons_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // buttons_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> buttons_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> buttons_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> buttons_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> buttons_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> buttons_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // buttons_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // buttons_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> buttons_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] buttons_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // buttons_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> buttons_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // buttons_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> buttons_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // solenoid_out_s1_translator:uav_waitrequest -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> solenoid_out_s1_translator:uav_burstcount
	wire   [31:0] solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> solenoid_out_s1_translator:uav_writedata
	wire   [26:0] solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_address -> solenoid_out_s1_translator:uav_address
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_write -> solenoid_out_s1_translator:uav_write
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_lock -> solenoid_out_s1_translator:uav_lock
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_read -> solenoid_out_s1_translator:uav_read
	wire   [31:0] solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // solenoid_out_s1_translator:uav_readdata -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // solenoid_out_s1_translator:uav_readdatavalid -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> solenoid_out_s1_translator:uav_debugaccess
	wire    [3:0] solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // solenoid_out_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> solenoid_out_s1_translator:uav_byteenable
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [104:0] solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [104:0] solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] solenoid_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // pwm_generator_0_avalon_slave_control_translator:uav_waitrequest -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_burstcount;              // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_burstcount -> pwm_generator_0_avalon_slave_control_translator:uav_burstcount
	wire    [7:0] pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_writedata;               // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_writedata -> pwm_generator_0_avalon_slave_control_translator:uav_writedata
	wire   [26:0] pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_address;                 // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_address -> pwm_generator_0_avalon_slave_control_translator:uav_address
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_write;                   // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_write -> pwm_generator_0_avalon_slave_control_translator:uav_write
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_lock;                    // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_lock -> pwm_generator_0_avalon_slave_control_translator:uav_lock
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_read;                    // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_read -> pwm_generator_0_avalon_slave_control_translator:uav_read
	wire    [7:0] pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_readdata;                // pwm_generator_0_avalon_slave_control_translator:uav_readdata -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // pwm_generator_0_avalon_slave_control_translator:uav_readdatavalid -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pwm_generator_0_avalon_slave_control_translator:uav_debugaccess
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_byteenable;              // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:m0_byteenable -> pwm_generator_0_avalon_slave_control_translator:uav_byteenable
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_valid;            // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rf_source_valid -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [77:0] pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_data;             // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rf_source_data -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_ready;            // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [77:0] pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [7:0] pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // nios2_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                            // nios2_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // nios2_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [103:0] nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                             // nios2_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router:sink_ready -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                             // nios2_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                   // nios2_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                           // nios2_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [103:0] nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                    // nios2_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                   // addr_router_001:sink_ready -> nios2_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                              // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [103:0] nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                               // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router:sink_ready -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [103:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_001:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [85:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_002:sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [103:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_003:sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [103:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_004:sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                     // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [103:0] altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                                      // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_005:sink_ready -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [103:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_006:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [103:0] green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // green_leds_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_007:sink_ready -> green_leds_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // switch_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                              // switch_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // switch_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [103:0] switch_s1_translator_avalon_universal_slave_0_agent_rp_data;                                               // switch_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          switch_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_008:sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_valid;                               // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [103:0] de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_data;                                // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_009:sink_ready -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid;                             // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [103:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data;                              // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_010:sink_ready -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [103:0] timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_011:sink_ready -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_valid;                    // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [103:0] pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_data;                     // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_012:sink_ready -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_valid;                      // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [103:0] pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_data;                       // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_013:sink_ready -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:rp_ready
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // buttons_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                             // buttons_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // buttons_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [103:0] buttons_s1_translator_avalon_universal_slave_0_agent_rp_data;                                              // buttons_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          buttons_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router_014:sink_ready -> buttons_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [103:0] solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // solenoid_out_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_015:sink_ready -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_valid;                   // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire   [76:0] pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_data;                    // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_016:sink_ready -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                                         // burst_adapter:source0_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                               // burst_adapter:source0_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                       // burst_adapter:source0_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [85:0] burst_adapter_source0_data;                                                                                // burst_adapter:source0_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                               // sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [16:0] burst_adapter_source0_channel;                                                                             // burst_adapter:source0_channel -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                     // burst_adapter_001:source0_endofpacket -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                           // burst_adapter_001:source0_valid -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                   // burst_adapter_001:source0_startofpacket -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [76:0] burst_adapter_001_source0_data;                                                                            // burst_adapter_001:source0_data -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                           // pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [16:0] burst_adapter_001_source0_channel;                                                                         // burst_adapter_001:source0_channel -> pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                            // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, crosser:in_reset, crosser_001:out_reset, de0_nano_adc_0:reset, de0_nano_adc_0_adc_slave_translator:reset, de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:reset, de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, green_leds:reset_n, green_leds_s1_translator:reset, green_leds_s1_translator_avalon_universal_slave_0_agent:reset, green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_003:reset, id_router_004:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_0:reset_n, nios2_0_data_master_translator:reset, nios2_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_0_instruction_master_translator:reset, nios2_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_0_jtag_debug_module_translator:reset, nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, switch:reset_n, switch_s1_translator:reset, switch_s1_translator_avalon_universal_slave_0_agent:reset, switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sys_clk_timer:reset_n, sys_clk_timer_s1_translator:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_qsys_0:reset_n, sysid_qsys_0_control_slave_translator:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_001_reset_out_reset;                                                                        // rst_controller_001:reset_out -> [altpll_0:reset, altpll_0_pll_slave_translator:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_001:in_reset, id_router_005:reset, rsp_xbar_demux_005:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                           // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                 // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                         // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [103:0] cmd_xbar_demux_src0_data;                                                                                  // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [16:0] cmd_xbar_demux_src0_channel;                                                                               // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                 // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                           // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                 // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                         // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [103:0] cmd_xbar_demux_src1_data;                                                                                  // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [16:0] cmd_xbar_demux_src1_channel;                                                                               // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                 // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                           // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                 // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                         // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [103:0] cmd_xbar_demux_src2_data;                                                                                  // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [16:0] cmd_xbar_demux_src2_channel;                                                                               // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                 // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                       // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                             // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                     // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src0_data;                                                                              // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [16:0] cmd_xbar_demux_001_src0_channel;                                                                           // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                             // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                       // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                             // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                     // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src1_data;                                                                              // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [16:0] cmd_xbar_demux_001_src1_channel;                                                                           // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                             // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                       // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                             // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                     // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src2_data;                                                                              // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [16:0] cmd_xbar_demux_001_src2_channel;                                                                           // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                             // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                       // cmd_xbar_demux_001:src3_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                             // cmd_xbar_demux_001:src3_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                     // cmd_xbar_demux_001:src3_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src3_data;                                                                              // cmd_xbar_demux_001:src3_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src3_channel;                                                                           // cmd_xbar_demux_001:src3_channel -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                       // cmd_xbar_demux_001:src4_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                             // cmd_xbar_demux_001:src4_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                     // cmd_xbar_demux_001:src4_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src4_data;                                                                              // cmd_xbar_demux_001:src4_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src4_channel;                                                                           // cmd_xbar_demux_001:src4_channel -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                       // cmd_xbar_demux_001:src6_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                             // cmd_xbar_demux_001:src6_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                     // cmd_xbar_demux_001:src6_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src6_data;                                                                              // cmd_xbar_demux_001:src6_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src6_channel;                                                                           // cmd_xbar_demux_001:src6_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                       // cmd_xbar_demux_001:src7_endofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                             // cmd_xbar_demux_001:src7_valid -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                     // cmd_xbar_demux_001:src7_startofpacket -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src7_data;                                                                              // cmd_xbar_demux_001:src7_data -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src7_channel;                                                                           // cmd_xbar_demux_001:src7_channel -> green_leds_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                       // cmd_xbar_demux_001:src8_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                             // cmd_xbar_demux_001:src8_valid -> switch_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                     // cmd_xbar_demux_001:src8_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src8_data;                                                                              // cmd_xbar_demux_001:src8_data -> switch_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src8_channel;                                                                           // cmd_xbar_demux_001:src8_channel -> switch_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                       // cmd_xbar_demux_001:src9_endofpacket -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                             // cmd_xbar_demux_001:src9_valid -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                     // cmd_xbar_demux_001:src9_startofpacket -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src9_data;                                                                              // cmd_xbar_demux_001:src9_data -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src9_channel;                                                                           // cmd_xbar_demux_001:src9_channel -> de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                      // cmd_xbar_demux_001:src10_endofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                            // cmd_xbar_demux_001:src10_valid -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                    // cmd_xbar_demux_001:src10_startofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src10_data;                                                                             // cmd_xbar_demux_001:src10_data -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src10_channel;                                                                          // cmd_xbar_demux_001:src10_channel -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                      // cmd_xbar_demux_001:src11_endofpacket -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                            // cmd_xbar_demux_001:src11_valid -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                    // cmd_xbar_demux_001:src11_startofpacket -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src11_data;                                                                             // cmd_xbar_demux_001:src11_data -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src11_channel;                                                                          // cmd_xbar_demux_001:src11_channel -> timestamp_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                      // cmd_xbar_demux_001:src12_endofpacket -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                            // cmd_xbar_demux_001:src12_valid -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                    // cmd_xbar_demux_001:src12_startofpacket -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src12_data;                                                                             // cmd_xbar_demux_001:src12_data -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src12_channel;                                                                          // cmd_xbar_demux_001:src12_channel -> pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                                      // cmd_xbar_demux_001:src13_endofpacket -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                            // cmd_xbar_demux_001:src13_valid -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                                    // cmd_xbar_demux_001:src13_startofpacket -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src13_data;                                                                             // cmd_xbar_demux_001:src13_data -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src13_channel;                                                                          // cmd_xbar_demux_001:src13_channel -> pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                                      // cmd_xbar_demux_001:src14_endofpacket -> buttons_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                            // cmd_xbar_demux_001:src14_valid -> buttons_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                                    // cmd_xbar_demux_001:src14_startofpacket -> buttons_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src14_data;                                                                             // cmd_xbar_demux_001:src14_data -> buttons_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src14_channel;                                                                          // cmd_xbar_demux_001:src14_channel -> buttons_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                                      // cmd_xbar_demux_001:src15_endofpacket -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                            // cmd_xbar_demux_001:src15_valid -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                                    // cmd_xbar_demux_001:src15_startofpacket -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src15_data;                                                                             // cmd_xbar_demux_001:src15_data -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_demux_001_src15_channel;                                                                          // cmd_xbar_demux_001:src15_channel -> solenoid_out_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                                      // cmd_xbar_demux_001:src16_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                            // cmd_xbar_demux_001:src16_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                                    // cmd_xbar_demux_001:src16_startofpacket -> width_adapter_002:in_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src16_data;                                                                             // cmd_xbar_demux_001:src16_data -> width_adapter_002:in_data
	wire   [16:0] cmd_xbar_demux_001_src16_channel;                                                                          // cmd_xbar_demux_001:src16_channel -> width_adapter_002:in_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                           // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                 // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                         // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [103:0] rsp_xbar_demux_src0_data;                                                                                  // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [16:0] rsp_xbar_demux_src0_channel;                                                                               // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                 // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                           // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                 // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                         // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [103:0] rsp_xbar_demux_src1_data;                                                                                  // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [16:0] rsp_xbar_demux_src1_channel;                                                                               // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                 // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                       // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                             // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                     // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [103:0] rsp_xbar_demux_001_src0_data;                                                                              // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [16:0] rsp_xbar_demux_001_src0_channel;                                                                           // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                             // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                       // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                             // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                     // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [103:0] rsp_xbar_demux_001_src1_data;                                                                              // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [16:0] rsp_xbar_demux_001_src1_channel;                                                                           // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                             // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                       // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                             // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                     // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [103:0] rsp_xbar_demux_002_src0_data;                                                                              // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [16:0] rsp_xbar_demux_002_src0_channel;                                                                           // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                             // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                       // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                             // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                     // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [103:0] rsp_xbar_demux_002_src1_data;                                                                              // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [16:0] rsp_xbar_demux_002_src1_channel;                                                                           // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                             // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                       // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                             // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                     // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [103:0] rsp_xbar_demux_003_src0_data;                                                                              // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [16:0] rsp_xbar_demux_003_src0_channel;                                                                           // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                             // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                       // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                             // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                     // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [103:0] rsp_xbar_demux_004_src0_data;                                                                              // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [16:0] rsp_xbar_demux_004_src0_channel;                                                                           // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                             // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                       // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                             // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                     // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [103:0] rsp_xbar_demux_006_src0_data;                                                                              // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [16:0] rsp_xbar_demux_006_src0_channel;                                                                           // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                             // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                       // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                             // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                     // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [103:0] rsp_xbar_demux_007_src0_data;                                                                              // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [16:0] rsp_xbar_demux_007_src0_channel;                                                                           // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                             // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                       // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                             // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                     // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [103:0] rsp_xbar_demux_008_src0_data;                                                                              // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [16:0] rsp_xbar_demux_008_src0_channel;                                                                           // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                             // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                       // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                             // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                     // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [103:0] rsp_xbar_demux_009_src0_data;                                                                              // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [16:0] rsp_xbar_demux_009_src0_channel;                                                                           // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                             // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                       // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                             // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                     // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [103:0] rsp_xbar_demux_010_src0_data;                                                                              // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [16:0] rsp_xbar_demux_010_src0_channel;                                                                           // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                             // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                       // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                             // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                     // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [103:0] rsp_xbar_demux_011_src0_data;                                                                              // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [16:0] rsp_xbar_demux_011_src0_channel;                                                                           // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                             // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                       // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                             // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                     // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [103:0] rsp_xbar_demux_012_src0_data;                                                                              // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [16:0] rsp_xbar_demux_012_src0_channel;                                                                           // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                             // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                       // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                             // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                     // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [103:0] rsp_xbar_demux_013_src0_data;                                                                              // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire   [16:0] rsp_xbar_demux_013_src0_channel;                                                                           // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                             // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                       // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                             // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                     // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [103:0] rsp_xbar_demux_014_src0_data;                                                                              // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire   [16:0] rsp_xbar_demux_014_src0_channel;                                                                           // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                             // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                       // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                             // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                     // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [103:0] rsp_xbar_demux_015_src0_data;                                                                              // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire   [16:0] rsp_xbar_demux_015_src0_channel;                                                                           // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                             // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                       // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                             // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                     // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [103:0] rsp_xbar_demux_016_src0_data;                                                                              // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire   [16:0] rsp_xbar_demux_016_src0_channel;                                                                           // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                             // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          addr_router_src_endofpacket;                                                                               // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                                     // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                             // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [103:0] addr_router_src_data;                                                                                      // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [16:0] addr_router_src_channel;                                                                                   // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                                     // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                              // rsp_xbar_mux:src_endofpacket -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                    // rsp_xbar_mux:src_valid -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                            // rsp_xbar_mux:src_startofpacket -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [103:0] rsp_xbar_mux_src_data;                                                                                     // rsp_xbar_mux:src_data -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [16:0] rsp_xbar_mux_src_channel;                                                                                  // rsp_xbar_mux:src_channel -> nios2_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                                    // nios2_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                           // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                 // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                         // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [103:0] addr_router_001_src_data;                                                                                  // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [16:0] addr_router_001_src_channel;                                                                               // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                 // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                          // rsp_xbar_mux_001:src_endofpacket -> nios2_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                // rsp_xbar_mux_001:src_valid -> nios2_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                        // rsp_xbar_mux_001:src_startofpacket -> nios2_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [103:0] rsp_xbar_mux_001_src_data;                                                                                 // rsp_xbar_mux_001:src_data -> nios2_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [16:0] rsp_xbar_mux_001_src_channel;                                                                              // rsp_xbar_mux_001:src_channel -> nios2_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                // nios2_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                              // cmd_xbar_mux:src_endofpacket -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                    // cmd_xbar_mux:src_valid -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                            // cmd_xbar_mux:src_startofpacket -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_mux_src_data;                                                                                     // cmd_xbar_mux:src_data -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_mux_src_channel;                                                                                  // cmd_xbar_mux:src_channel -> nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                    // nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                 // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                       // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                               // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [103:0] id_router_src_data;                                                                                        // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [16:0] id_router_src_channel;                                                                                     // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                       // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                          // cmd_xbar_mux_001:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                // cmd_xbar_mux_001:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                        // cmd_xbar_mux_001:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] cmd_xbar_mux_001_src_data;                                                                                 // cmd_xbar_mux_001:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] cmd_xbar_mux_001_src_channel;                                                                              // cmd_xbar_mux_001:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                             // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                   // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                           // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [103:0] id_router_001_src_data;                                                                                    // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [16:0] id_router_001_src_channel;                                                                                 // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                   // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_003_src_endofpacket;                                                                             // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                   // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                           // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [103:0] id_router_003_src_data;                                                                                    // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [16:0] id_router_003_src_channel;                                                                                 // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                   // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                             // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                   // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                           // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [103:0] id_router_004_src_data;                                                                                    // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [16:0] id_router_004_src_channel;                                                                                 // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                   // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          crosser_out_ready;                                                                                         // altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_005_src_endofpacket;                                                                             // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                   // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                           // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [103:0] id_router_005_src_data;                                                                                    // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [16:0] id_router_005_src_channel;                                                                                 // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                   // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                             // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                   // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                           // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [103:0] id_router_006_src_data;                                                                                    // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [16:0] id_router_006_src_channel;                                                                                 // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                   // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                             // green_leds_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                             // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                   // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                           // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [103:0] id_router_007_src_data;                                                                                    // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [16:0] id_router_007_src_channel;                                                                                 // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                   // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                             // switch_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                             // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                   // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                           // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [103:0] id_router_008_src_data;                                                                                    // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [16:0] id_router_008_src_channel;                                                                                 // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                   // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                             // de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_009_src_endofpacket;                                                                             // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                   // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                           // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [103:0] id_router_009_src_data;                                                                                    // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [16:0] id_router_009_src_channel;                                                                                 // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                   // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src10_ready;                                                                            // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire          id_router_010_src_endofpacket;                                                                             // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                   // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                           // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [103:0] id_router_010_src_data;                                                                                    // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [16:0] id_router_010_src_channel;                                                                                 // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                   // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_001_src11_ready;                                                                            // timestamp_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire          id_router_011_src_endofpacket;                                                                             // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                   // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                           // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [103:0] id_router_011_src_data;                                                                                    // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [16:0] id_router_011_src_channel;                                                                                 // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                   // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                            // pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                             // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                   // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                           // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [103:0] id_router_012_src_data;                                                                                    // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [16:0] id_router_012_src_channel;                                                                                 // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                   // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_001_src13_ready;                                                                            // pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire          id_router_013_src_endofpacket;                                                                             // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                   // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                           // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [103:0] id_router_013_src_data;                                                                                    // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [16:0] id_router_013_src_channel;                                                                                 // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                   // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_001_src14_ready;                                                                            // buttons_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire          id_router_014_src_endofpacket;                                                                             // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                   // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                           // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [103:0] id_router_014_src_data;                                                                                    // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [16:0] id_router_014_src_channel;                                                                                 // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                   // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_001_src15_ready;                                                                            // solenoid_out_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	wire          id_router_015_src_endofpacket;                                                                             // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                   // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                           // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [103:0] id_router_015_src_data;                                                                                    // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [16:0] id_router_015_src_channel;                                                                                 // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                   // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                          // cmd_xbar_mux_002:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                // cmd_xbar_mux_002:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                        // cmd_xbar_mux_002:src_startofpacket -> width_adapter:in_startofpacket
	wire  [103:0] cmd_xbar_mux_002_src_data;                                                                                 // cmd_xbar_mux_002:src_data -> width_adapter:in_data
	wire   [16:0] cmd_xbar_mux_002_src_channel;                                                                              // cmd_xbar_mux_002:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                // width_adapter:in_ready -> cmd_xbar_mux_002:src_ready
	wire          width_adapter_src_endofpacket;                                                                             // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                   // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                           // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [85:0] width_adapter_src_data;                                                                                    // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                                   // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [16:0] width_adapter_src_channel;                                                                                 // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_002_src_endofpacket;                                                                             // id_router_002:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_002_src_valid;                                                                                   // id_router_002:src_valid -> width_adapter_001:in_valid
	wire          id_router_002_src_startofpacket;                                                                           // id_router_002:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [85:0] id_router_002_src_data;                                                                                    // id_router_002:src_data -> width_adapter_001:in_data
	wire   [16:0] id_router_002_src_channel;                                                                                 // id_router_002:src_channel -> width_adapter_001:in_channel
	wire          id_router_002_src_ready;                                                                                   // width_adapter_001:in_ready -> id_router_002:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                         // width_adapter_001:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                               // width_adapter_001:out_valid -> rsp_xbar_demux_002:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                       // width_adapter_001:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [103:0] width_adapter_001_src_data;                                                                                // width_adapter_001:out_data -> rsp_xbar_demux_002:sink_data
	wire          width_adapter_001_src_ready;                                                                               // rsp_xbar_demux_002:sink_ready -> width_adapter_001:out_ready
	wire   [16:0] width_adapter_001_src_channel;                                                                             // width_adapter_001:out_channel -> rsp_xbar_demux_002:sink_channel
	wire          cmd_xbar_demux_001_src16_ready;                                                                            // width_adapter_002:in_ready -> cmd_xbar_demux_001:src16_ready
	wire          width_adapter_002_src_endofpacket;                                                                         // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                               // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                       // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [76:0] width_adapter_002_src_data;                                                                                // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire          width_adapter_002_src_ready;                                                                               // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire   [16:0] width_adapter_002_src_channel;                                                                             // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          id_router_016_src_endofpacket;                                                                             // id_router_016:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_016_src_valid;                                                                                   // id_router_016:src_valid -> width_adapter_003:in_valid
	wire          id_router_016_src_startofpacket;                                                                           // id_router_016:src_startofpacket -> width_adapter_003:in_startofpacket
	wire   [76:0] id_router_016_src_data;                                                                                    // id_router_016:src_data -> width_adapter_003:in_data
	wire   [16:0] id_router_016_src_channel;                                                                                 // id_router_016:src_channel -> width_adapter_003:in_channel
	wire          id_router_016_src_ready;                                                                                   // width_adapter_003:in_ready -> id_router_016:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                         // width_adapter_003:out_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                               // width_adapter_003:out_valid -> rsp_xbar_demux_016:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                                       // width_adapter_003:out_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [103:0] width_adapter_003_src_data;                                                                                // width_adapter_003:out_data -> rsp_xbar_demux_016:sink_data
	wire          width_adapter_003_src_ready;                                                                               // rsp_xbar_demux_016:sink_ready -> width_adapter_003:out_ready
	wire   [16:0] width_adapter_003_src_channel;                                                                             // width_adapter_003:out_channel -> rsp_xbar_demux_016:sink_channel
	wire          crosser_out_endofpacket;                                                                                   // crosser:out_endofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                         // crosser:out_valid -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                                 // crosser:out_startofpacket -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [103:0] crosser_out_data;                                                                                          // crosser:out_data -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [16:0] crosser_out_channel;                                                                                       // crosser:out_channel -> altpll_0_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                       // cmd_xbar_demux_001:src5_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                             // cmd_xbar_demux_001:src5_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                     // cmd_xbar_demux_001:src5_startofpacket -> crosser:in_startofpacket
	wire  [103:0] cmd_xbar_demux_001_src5_data;                                                                              // cmd_xbar_demux_001:src5_data -> crosser:in_data
	wire   [16:0] cmd_xbar_demux_001_src5_channel;                                                                           // cmd_xbar_demux_001:src5_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src5_ready;                                                                             // crosser:in_ready -> cmd_xbar_demux_001:src5_ready
	wire          crosser_001_out_endofpacket;                                                                               // crosser_001:out_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          crosser_001_out_valid;                                                                                     // crosser_001:out_valid -> rsp_xbar_mux_001:sink5_valid
	wire          crosser_001_out_startofpacket;                                                                             // crosser_001:out_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [103:0] crosser_001_out_data;                                                                                      // crosser_001:out_data -> rsp_xbar_mux_001:sink5_data
	wire   [16:0] crosser_001_out_channel;                                                                                   // crosser_001:out_channel -> rsp_xbar_mux_001:sink5_channel
	wire          crosser_001_out_ready;                                                                                     // rsp_xbar_mux_001:sink5_ready -> crosser_001:out_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                       // rsp_xbar_demux_005:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                             // rsp_xbar_demux_005:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                     // rsp_xbar_demux_005:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [103:0] rsp_xbar_demux_005_src0_data;                                                                              // rsp_xbar_demux_005:src0_data -> crosser_001:in_data
	wire   [16:0] rsp_xbar_demux_005_src0_channel;                                                                           // rsp_xbar_demux_005:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                             // crosser_001:in_ready -> rsp_xbar_demux_005:src0_ready
	wire          irq_mapper_receiver0_irq;                                                                                  // sys_clk_timer:irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                  // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                  // rs232_0:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                  // timestamp_timer:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                                  // buttons:irq -> irq_mapper:receiver4_irq
	wire   [31:0] nios2_0_d_irq_irq;                                                                                         // irq_mapper:sender_irq -> nios2_0:d_irq

	niosII_system_nios2_0 nios2_0 (
		.clk                                   (altpll_0_c1_clk),                                                        //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                        //                   reset_n.reset_n
		.d_address                             (nios2_0_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_0_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_0_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_0_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_0_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_0_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_0_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_0_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_0_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_0_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_0_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_0_instruction_master_waitrequest),                                 //                          .waitrequest
		.d_irq                                 (nios2_0_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_0_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                        // custom_instruction_master.readra
	);

	niosII_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c1_clk),                                               //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                                 // reset1.reset
	);

	niosII_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c1_clk),                                                    //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                                    //         reset.reset_n
		.readdata (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	niosII_system_sys_clk_timer sys_clk_timer (
		.clk        (altpll_0_c1_clk),                                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                            // reset.reset_n
		.address    (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~sys_clk_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                                    //   irq.irq
	);

	niosII_system_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c1_clk),                                                          //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                                  //               irq.irq
	);

	niosII_system_green_leds green_leds (
		.clk        (altpll_0_c1_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (green_leds_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~green_leds_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (green_leds_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (green_leds_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (green_leds_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_green_leds)                             // external_connection.export
	);

	niosII_system_switch switch (
		.clk      (altpll_0_c1_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (switch_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (switch_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (in_port_to_the_switch)                              // external_connection.export
	);

	niosII_system_altpll_0 altpll_0 (
		.clk       (clk_0),                                                       //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),                          // inclk_interface_reset.reset
		.read      (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (altpll_0_c0_out),                                             //                    c0.clk
		.c1        (altpll_0_c1_clk),                                             //                    c1.clk
		.areset    (areset_to_the_altpll_0),                                      //        areset_conduit.export
		.locked    (locked_from_the_altpll_0),                                    //        locked_conduit.export
		.phasedone (phasedone_from_the_altpll_0)                                  //     phasedone_conduit.export
	);

	niosII_system_de0_nano_adc_0 de0_nano_adc_0 (
		.clock       (altpll_0_c1_clk),                                                     //                clk.clk
		.reset       (rst_controller_reset_out_reset),                                      //              reset.reset
		.write       (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_write),       //          adc_slave.write
		.readdata    (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.writedata   (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.address     (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_address),     //                   .address
		.waitrequest (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.read        (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.adc_sclk    (adc_sclk_from_the_de0_nano_adc_0),                                    // external_interface.export
		.adc_cs_n    (adc_cs_n_from_the_de0_nano_adc_0),                                    //                   .export
		.adc_dout    (adc_dout_to_the_de0_nano_adc_0),                                      //                   .export
		.adc_din     (adc_din_from_the_de0_nano_adc_0)                                      //                   .export
	);

	niosII_system_sdram_0 sdram_0 (
		.clk            (altpll_0_c1_clk),                                         //   clk.clk
		.reset_n        (~nios2_0_jtag_debug_module_reset_reset),                  // reset.reset_n
		.az_addr        (sdram_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_0_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_0_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_0_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_0_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_0_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_0_wire_dq),                                         //      .export
		.zs_dqm         (sdram_0_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_0_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_0_wire_we_n)                                        //      .export
	);

	niosII_system_rs232_0 rs232_0 (
		.clk        (altpll_0_c1_clk),                                                      //        clock_reset.clk
		.reset      (nios2_0_jtag_debug_module_reset_reset),                                //  clock_reset_reset.reset
		.address    (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_address),    // avalon_rs232_slave.address
		.chipselect (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.byteenable (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable), //                   .byteenable
		.read       (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write      (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata  (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata   (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver2_irq),                                             //          interrupt.irq
		.UART_RXD   (rs232_0_external_interface_RXD),                                       // external_interface.export
		.UART_TXD   (rs232_0_external_interface_TXD)                                        //                   .export
	);

	niosII_system_timestamp_timer timestamp_timer (
		.clk        (altpll_0_c1_clk),                                              //   clk.clk
		.reset_n    (~nios2_0_jtag_debug_module_reset_reset),                       // reset.reset_n
		.address    (timestamp_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timestamp_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timestamp_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timestamp_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timestamp_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                                      //   irq.irq
	);

	pwm_generator pwm_generator_0 (
		.reset            (nios2_0_jtag_debug_module_reset_reset),                                         //                reset.reset
		.clock            (altpll_0_c1_clk),                                                               //           clock_sink.clk
		.pwm_out          (pwm_generator_0_pwm_out_export),                                                //              pwm_out.export
		.write_en_period  (pwm_generator_0_avalon_slave_period_translator_avalon_anti_slave_0_write),      //  avalon_slave_period.write
		.period_in        (pwm_generator_0_avalon_slave_period_translator_avalon_anti_slave_0_writedata),  //                     .writedata
		.write_en_duty    (pwm_generator_0_avalon_slave_duty_translator_avalon_anti_slave_0_write),        //    avalon_slave_duty.write
		.duty_in          (pwm_generator_0_avalon_slave_duty_translator_avalon_anti_slave_0_writedata),    //                     .writedata
		.write_en_control (pwm_generator_0_avalon_slave_control_translator_avalon_anti_slave_0_write),     // avalon_slave_control.write
		.control_in       (pwm_generator_0_avalon_slave_control_translator_avalon_anti_slave_0_writedata)  //                     .writedata
	);

	niosII_system_buttons buttons (
		.clk        (altpll_0_c1_clk),                                      //                 clk.clk
		.reset_n    (~nios2_0_jtag_debug_module_reset_reset),               //               reset.reset_n
		.address    (buttons_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~buttons_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (buttons_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (buttons_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (buttons_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (buttons_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                              //                 irq.irq
	);

	niosII_system_solenoid_out solenoid_out (
		.clk        (altpll_0_c1_clk),                                           //                 clk.clk
		.reset_n    (~nios2_0_jtag_debug_module_reset_reset),                    //               reset.reset_n
		.address    (solenoid_out_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~solenoid_out_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (solenoid_out_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (solenoid_out_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (solenoid_out_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (solenoid_out_external_connection_export)                    // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (27),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_0_instruction_master_translator (
		.clk                   (altpll_0_c1_clk),                                                               //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                //                     reset.reset
		.uav_address           (nios2_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_0_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount         (1'b1),                                                                          //               (terminated)
		.av_byteenable         (4'b1111),                                                                       //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                          //               (terminated)
		.av_begintransfer      (1'b0),                                                                          //               (terminated)
		.av_chipselect         (1'b0),                                                                          //               (terminated)
		.av_readdatavalid      (),                                                                              //               (terminated)
		.av_write              (1'b0),                                                                          //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                          //               (terminated)
		.av_lock               (1'b0),                                                                          //               (terminated)
		.av_debugaccess        (1'b0),                                                                          //               (terminated)
		.uav_clken             (),                                                                              //               (terminated)
		.av_clken              (1'b1)                                                                           //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (27),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2_0_data_master_translator (
		.clk                   (altpll_0_c1_clk),                                                        //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                     reset.reset
		.uav_address           (nios2_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_0_data_master_read),                                               //                          .read
		.av_readdata           (nios2_0_data_master_readdata),                                           //                          .readdata
		.av_write              (nios2_0_data_master_write),                                              //                          .write
		.av_writedata          (nios2_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                   //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                   //               (terminated)
		.av_begintransfer      (1'b0),                                                                   //               (terminated)
		.av_chipselect         (1'b0),                                                                   //               (terminated)
		.av_readdatavalid      (),                                                                       //               (terminated)
		.av_lock               (1'b0),                                                                   //               (terminated)
		.uav_clken             (),                                                                       //               (terminated)
		.av_clken              (1'b1)                                                                    //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_0_jtag_debug_module_translator (
		.clk                   (altpll_0_c1_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_0_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                       //                      clk.clk
		.reset                 (nios2_0_jtag_debug_module_reset_reset),                                 //                    reset.reset
		.uav_address           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_0_control_slave_translator (
		.clk                   (altpll_0_c1_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                                      //              (terminated)
		.av_read               (),                                                                                      //              (terminated)
		.av_writedata          (),                                                                                      //              (terminated)
		.av_begintransfer      (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_byteenable         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_chipselect         (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sys_clk_timer_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sys_clk_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_byteenable         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.av_clken              (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altpll_0_pll_slave_translator (
		.clk                   (clk_0),                                                                         //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                            //                    reset.reset
		.uav_address           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (altpll_0_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (altpll_0_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (altpll_0_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (altpll_0_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (altpll_0_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_chipselect         (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (altpll_0_c1_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) green_leds_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (green_leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (green_leds_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (green_leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (green_leds_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (green_leds_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (switch_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (switch_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (switch_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (switch_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (switch_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (switch_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_writedata          (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) de0_nano_adc_0_adc_slave_translator (
		.clk                   (altpll_0_c1_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (de0_nano_adc_0_adc_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_byteenable         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_chipselect         (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rs232_0_avalon_rs232_slave_translator (
		.clk                   (altpll_0_c1_clk),                                                                       //                      clk.clk
		.reset                 (nios2_0_jtag_debug_module_reset_reset),                                                 //                    reset.reset
		.uav_address           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timestamp_timer_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                               //                      clk.clk
		.reset                 (nios2_0_jtag_debug_module_reset_reset),                                         //                    reset.reset
		.uav_address           (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timestamp_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timestamp_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timestamp_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timestamp_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timestamp_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                              //              (terminated)
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_byteenable         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_waitrequest        (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pwm_generator_0_avalon_slave_period_translator (
		.clk                   (altpll_0_c1_clk),                                                                                //                      clk.clk
		.reset                 (nios2_0_jtag_debug_module_reset_reset),                                                          //                    reset.reset
		.uav_address           (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (pwm_generator_0_avalon_slave_period_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (pwm_generator_0_avalon_slave_period_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_address            (),                                                                                               //              (terminated)
		.av_read               (),                                                                                               //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                                           //              (terminated)
		.av_begintransfer      (),                                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                                               //              (terminated)
		.av_burstcount         (),                                                                                               //              (terminated)
		.av_byteenable         (),                                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                                               //              (terminated)
		.av_lock               (),                                                                                               //              (terminated)
		.av_chipselect         (),                                                                                               //              (terminated)
		.av_clken              (),                                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                                           //              (terminated)
		.av_debugaccess        (),                                                                                               //              (terminated)
		.av_outputenable       ()                                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pwm_generator_0_avalon_slave_duty_translator (
		.clk                   (altpll_0_c1_clk),                                                                              //                      clk.clk
		.reset                 (nios2_0_jtag_debug_module_reset_reset),                                                        //                    reset.reset
		.uav_address           (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (pwm_generator_0_avalon_slave_duty_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (pwm_generator_0_avalon_slave_duty_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_address            (),                                                                                             //              (terminated)
		.av_read               (),                                                                                             //              (terminated)
		.av_readdata           (32'b11011110101011011101111010101101),                                                         //              (terminated)
		.av_begintransfer      (),                                                                                             //              (terminated)
		.av_beginbursttransfer (),                                                                                             //              (terminated)
		.av_burstcount         (),                                                                                             //              (terminated)
		.av_byteenable         (),                                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                                             //              (terminated)
		.av_lock               (),                                                                                             //              (terminated)
		.av_chipselect         (),                                                                                             //              (terminated)
		.av_clken              (),                                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                                         //              (terminated)
		.av_debugaccess        (),                                                                                             //              (terminated)
		.av_outputenable       ()                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) buttons_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                       //                      clk.clk
		.reset                 (nios2_0_jtag_debug_module_reset_reset),                                 //                    reset.reset
		.uav_address           (buttons_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (buttons_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (buttons_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (buttons_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (buttons_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (buttons_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (buttons_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (buttons_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (buttons_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (buttons_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (buttons_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (buttons_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (buttons_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (buttons_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (buttons_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (buttons_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) solenoid_out_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                            //                      clk.clk
		.reset                 (nios2_0_jtag_debug_module_reset_reset),                                      //                    reset.reset
		.uav_address           (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (solenoid_out_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (solenoid_out_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (solenoid_out_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (solenoid_out_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (solenoid_out_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                           //              (terminated)
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_burstcount         (),                                                                           //              (terminated)
		.av_byteenable         (),                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                       //              (terminated)
		.av_waitrequest        (1'b0),                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pwm_generator_0_avalon_slave_control_translator (
		.clk                   (altpll_0_c1_clk),                                                                                 //                      clk.clk
		.reset                 (nios2_0_jtag_debug_module_reset_reset),                                                           //                    reset.reset
		.uav_address           (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_write              (pwm_generator_0_avalon_slave_control_translator_avalon_anti_slave_0_write),                       //      avalon_anti_slave_0.write
		.av_writedata          (pwm_generator_0_avalon_slave_control_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_address            (),                                                                                                //              (terminated)
		.av_read               (),                                                                                                //              (terminated)
		.av_readdata           (8'b10101101),                                                                                     //              (terminated)
		.av_begintransfer      (),                                                                                                //              (terminated)
		.av_beginbursttransfer (),                                                                                                //              (terminated)
		.av_burstcount         (),                                                                                                //              (terminated)
		.av_byteenable         (),                                                                                                //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                            //              (terminated)
		.av_waitrequest        (1'b0),                                                                                            //              (terminated)
		.av_writebyteenable    (),                                                                                                //              (terminated)
		.av_lock               (),                                                                                                //              (terminated)
		.av_chipselect         (),                                                                                                //              (terminated)
		.av_clken              (),                                                                                                //              (terminated)
		.uav_clken             (1'b0),                                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                                //              (terminated)
		.av_outputenable       ()                                                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_BEGIN_BURST           (82),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.PKT_BURST_TYPE_H          (79),
		.PKT_BURST_TYPE_L          (78),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_TRANS_EXCLUSIVE       (68),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_THREAD_ID_H           (94),
		.PKT_THREAD_ID_L           (94),
		.PKT_CACHE_H               (101),
		.PKT_CACHE_L               (98),
		.PKT_DATA_SIDEBAND_H       (81),
		.PKT_DATA_SIDEBAND_L       (81),
		.PKT_QOS_H                 (83),
		.PKT_QOS_L                 (83),
		.PKT_ADDR_SIDEBAND_H       (80),
		.PKT_ADDR_SIDEBAND_L       (80),
		.ST_DATA_W                 (104),
		.ST_CHANNEL_W              (17),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) nios2_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c1_clk),                                                                        //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.av_address       (nios2_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_src_valid),                                                                 //        rp.valid
		.rp_data          (rsp_xbar_mux_src_data),                                                                  //          .data
		.rp_channel       (rsp_xbar_mux_src_channel),                                                               //          .channel
		.rp_startofpacket (rsp_xbar_mux_src_startofpacket),                                                         //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_src_endofpacket),                                                           //          .endofpacket
		.rp_ready         (rsp_xbar_mux_src_ready)                                                                  //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_BEGIN_BURST           (82),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.PKT_BURST_TYPE_H          (79),
		.PKT_BURST_TYPE_L          (78),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_TRANS_EXCLUSIVE       (68),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_THREAD_ID_H           (94),
		.PKT_THREAD_ID_L           (94),
		.PKT_CACHE_H               (101),
		.PKT_CACHE_L               (98),
		.PKT_DATA_SIDEBAND_H       (81),
		.PKT_DATA_SIDEBAND_L       (81),
		.PKT_QOS_H                 (83),
		.PKT_QOS_L                 (83),
		.PKT_ADDR_SIDEBAND_H       (80),
		.PKT_ADDR_SIDEBAND_L       (80),
		.ST_DATA_W                 (104),
		.ST_CHANNEL_W              (17),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) nios2_0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c1_clk),                                                                 //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.av_address       (nios2_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                      //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                       //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                    //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                              //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                                //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                       //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                       //                .channel
		.rf_sink_ready           (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                             //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (75),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (79),
		.PKT_PROTECTION_L          (77),
		.PKT_RESPONSE_STATUS_H     (85),
		.PKT_RESPONSE_STATUS_L     (84),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (86),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                 //             clk.clk
		.reset                   (nios2_0_jtag_debug_module_reset_reset),                                           //       clk_reset.reset
		.m0_address              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                     //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                     //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                      //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                               //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                   //                .channel
		.rf_sink_ready           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (87),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                 //       clk.clk
		.reset             (nios2_0_jtag_debug_module_reset_reset),                                           // clk_reset.reset
		.in_data           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                 //                .channel
		.rf_sink_ready           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                       //                .channel
		.rf_sink_ready           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_0),                                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                       //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                       //                .valid
		.cp_data                 (crosser_out_data),                                                                        //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                     //                .channel
		.rf_sink_ready           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_0),                                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_0),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                // clk_reset.reset
		.in_data           (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_startofpacket  (1'b0),                                                                              // (terminated)
		.in_endofpacket    (1'b0),                                                                              // (terminated)
		.out_startofpacket (),                                                                                  // (terminated)
		.out_endofpacket   (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) green_leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (green_leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                    //                .channel
		.rf_sink_ready           (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (green_leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (green_leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) switch_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (switch_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                //                .channel
		.rf_sink_ready           (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                                               //                .channel
		.rf_sink_ready           (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                 //             clk.clk
		.reset                   (nios2_0_jtag_debug_module_reset_reset),                                                           //       clk_reset.reset
		.m0_address              (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                                //                .channel
		.rf_sink_ready           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                 //       clk.clk
		.reset             (nios2_0_jtag_debug_module_reset_reset),                                                           // clk_reset.reset
		.in_data           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timestamp_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                         //             clk.clk
		.reset                   (nios2_0_jtag_debug_module_reset_reset),                                                   //       clk_reset.reset
		.m0_address              (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                        //                .channel
		.rf_sink_ready           (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                         //       clk.clk
		.reset             (nios2_0_jtag_debug_module_reset_reset),                                                   // clk_reset.reset
		.in_data           (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                          //             clk.clk
		.reset                   (nios2_0_jtag_debug_module_reset_reset),                                                                    //       clk_reset.reset
		.m0_address              (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                                           //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                                           //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                                            //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                                         //                .channel
		.rf_sink_ready           (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                          //       clk.clk
		.reset             (nios2_0_jtag_debug_module_reset_reset),                                                                    // clk_reset.reset
		.in_data           (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                                     // (terminated)
		.csr_readdata      (),                                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                     // (terminated)
		.almost_full_data  (),                                                                                                         // (terminated)
		.almost_empty_data (),                                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                                     // (terminated)
		.out_empty         (),                                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                                     // (terminated)
		.out_error         (),                                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                                     // (terminated)
		.out_channel       ()                                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                        //             clk.clk
		.reset                   (nios2_0_jtag_debug_module_reset_reset),                                                                  //       clk_reset.reset
		.m0_address              (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                                       //                .channel
		.rf_sink_ready           (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                        //       clk.clk
		.reset             (nios2_0_jtag_debug_module_reset_reset),                                                                  // clk_reset.reset
		.in_data           (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) buttons_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                 //             clk.clk
		.reset                   (nios2_0_jtag_debug_module_reset_reset),                                           //       clk_reset.reset
		.m0_address              (buttons_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (buttons_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (buttons_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (buttons_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (buttons_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (buttons_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (buttons_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (buttons_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (buttons_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (buttons_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (buttons_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (buttons_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (buttons_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (buttons_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (buttons_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (buttons_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                                //                .channel
		.rf_sink_ready           (buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (buttons_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (buttons_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (buttons_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (buttons_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (buttons_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (buttons_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                 //       clk.clk
		.reset             (nios2_0_jtag_debug_module_reset_reset),                                           // clk_reset.reset
		.in_data           (buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (buttons_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (buttons_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (82),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (84),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (74),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.PKT_BURST_SIZE_H          (77),
		.PKT_BURST_SIZE_L          (75),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (104),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) solenoid_out_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                      //             clk.clk
		.reset                   (nios2_0_jtag_debug_module_reset_reset),                                                //       clk_reset.reset
		.m0_address              (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (solenoid_out_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src15_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src15_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src15_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src15_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src15_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src15_channel),                                                     //                .channel
		.rf_sink_ready           (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (105),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                      //       clk.clk
		.reset             (nios2_0_jtag_debug_module_reset_reset),                                                // clk_reset.reset
		.in_data           (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (55),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (35),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (36),
		.PKT_TRANS_POSTED          (37),
		.PKT_TRANS_WRITE           (38),
		.PKT_TRANS_READ            (39),
		.PKT_TRANS_LOCK            (40),
		.PKT_SRC_ID_H              (61),
		.PKT_SRC_ID_L              (57),
		.PKT_DEST_ID_H             (66),
		.PKT_DEST_ID_L             (62),
		.PKT_BURSTWRAP_H           (47),
		.PKT_BURSTWRAP_L           (45),
		.PKT_BYTE_CNT_H            (44),
		.PKT_BYTE_CNT_L            (42),
		.PKT_PROTECTION_H          (70),
		.PKT_PROTECTION_L          (68),
		.PKT_RESPONSE_STATUS_H     (76),
		.PKT_RESPONSE_STATUS_L     (75),
		.PKT_BURST_SIZE_H          (50),
		.PKT_BURST_SIZE_L          (48),
		.ST_CHANNEL_W              (17),
		.ST_DATA_W                 (77),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                           //             clk.clk
		.reset                   (nios2_0_jtag_debug_module_reset_reset),                                                                     //       clk_reset.reset
		.m0_address              (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                                           //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                                           //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                            //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                                         //                .channel
		.rf_sink_ready           (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (78),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                           //       clk.clk
		.reset             (nios2_0_jtag_debug_module_reset_reset),                                                                     // clk_reset.reset
		.in_data           (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                                      // (terminated)
		.csr_readdata      (),                                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                      // (terminated)
		.almost_full_data  (),                                                                                                          // (terminated)
		.almost_empty_data (),                                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                                      // (terminated)
		.out_empty         (),                                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                                      // (terminated)
		.out_error         (),                                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                                      // (terminated)
		.out_channel       ()                                                                                                           // (terminated)
	);

	niosII_system_addr_router addr_router (
		.sink_ready         (nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                  //       src.ready
		.src_valid          (addr_router_src_valid),                                                                  //          .valid
		.src_data           (addr_router_src_data),                                                                   //          .data
		.src_channel        (addr_router_src_channel),                                                                //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                             //          .endofpacket
	);

	niosII_system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                       //          .valid
		.src_data           (addr_router_001_src_data),                                                        //          .data
		.src_channel        (addr_router_001_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                  //          .endofpacket
	);

	niosII_system_id_router id_router (
		.sink_ready         (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_src_valid),                                                                  //          .valid
		.src_data           (id_router_src_data),                                                                   //          .data
		.src_channel        (id_router_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                             //          .endofpacket
	);

	niosII_system_id_router id_router_001 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                        //       src.ready
		.src_valid          (id_router_001_src_valid),                                                        //          .valid
		.src_data           (id_router_001_src_data),                                                         //          .data
		.src_channel        (id_router_001_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                   //          .endofpacket
	);

	niosII_system_id_router_002 id_router_002 (
		.sink_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset),                                 // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                               //       src.ready
		.src_valid          (id_router_002_src_valid),                                               //          .valid
		.src_data           (id_router_002_src_data),                                                //          .data
		.src_channel        (id_router_002_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                          //          .endofpacket
	);

	niosII_system_id_router_003 id_router_003 (
		.sink_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                               //       src.ready
		.src_valid          (id_router_003_src_valid),                                                               //          .valid
		.src_data           (id_router_003_src_data),                                                                //          .data
		.src_channel        (id_router_003_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                          //          .endofpacket
	);

	niosII_system_id_router_003 id_router_004 (
		.sink_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                     //       src.ready
		.src_valid          (id_router_004_src_valid),                                                     //          .valid
		.src_data           (id_router_004_src_data),                                                      //          .data
		.src_channel        (id_router_004_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                //          .endofpacket
	);

	niosII_system_id_router_003 id_router_005 (
		.sink_ready         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altpll_0_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_0),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                       //       src.ready
		.src_valid          (id_router_005_src_valid),                                                       //          .valid
		.src_data           (id_router_005_src_data),                                                        //          .data
		.src_channel        (id_router_005_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                  //          .endofpacket
	);

	niosII_system_id_router_003 id_router_006 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                  //          .valid
		.src_data           (id_router_006_src_data),                                                                   //          .data
		.src_channel        (id_router_006_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                             //          .endofpacket
	);

	niosII_system_id_router_003 id_router_007 (
		.sink_ready         (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (green_leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                  //       src.ready
		.src_valid          (id_router_007_src_valid),                                                  //          .valid
		.src_data           (id_router_007_src_data),                                                   //          .data
		.src_channel        (id_router_007_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                             //          .endofpacket
	);

	niosII_system_id_router_003 id_router_008 (
		.sink_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                              //       src.ready
		.src_valid          (id_router_008_src_valid),                                              //          .valid
		.src_data           (id_router_008_src_data),                                               //          .data
		.src_channel        (id_router_008_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                         //          .endofpacket
	);

	niosII_system_id_router_003 id_router_009 (
		.sink_ready         (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (de0_nano_adc_0_adc_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                             //       src.ready
		.src_valid          (id_router_009_src_valid),                                                             //          .valid
		.src_data           (id_router_009_src_data),                                                              //          .data
		.src_channel        (id_router_009_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                        //          .endofpacket
	);

	niosII_system_id_router_003 id_router_010 (
		.sink_ready         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                                               //          .valid
		.src_data           (id_router_010_src_data),                                                                //          .data
		.src_channel        (id_router_010_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                          //          .endofpacket
	);

	niosII_system_id_router_003 id_router_011 (
		.sink_ready         (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timestamp_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                               //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset),                                         // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                       //       src.ready
		.src_valid          (id_router_011_src_valid),                                                       //          .valid
		.src_data           (id_router_011_src_data),                                                        //          .data
		.src_channel        (id_router_011_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                  //          .endofpacket
	);

	niosII_system_id_router_003 id_router_012 (
		.sink_ready         (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pwm_generator_0_avalon_slave_period_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                                //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                                        //       src.ready
		.src_valid          (id_router_012_src_valid),                                                                        //          .valid
		.src_data           (id_router_012_src_data),                                                                         //          .data
		.src_channel        (id_router_012_src_channel),                                                                      //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                                   //          .endofpacket
	);

	niosII_system_id_router_003 id_router_013 (
		.sink_ready         (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pwm_generator_0_avalon_slave_duty_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                              //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_013_src_valid),                                                                      //          .valid
		.src_data           (id_router_013_src_data),                                                                       //          .data
		.src_channel        (id_router_013_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                                 //          .endofpacket
	);

	niosII_system_id_router_003 id_router_014 (
		.sink_ready         (buttons_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (buttons_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (buttons_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (buttons_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (buttons_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset),                                 // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                               //       src.ready
		.src_valid          (id_router_014_src_valid),                                               //          .valid
		.src_data           (id_router_014_src_data),                                                //          .data
		.src_channel        (id_router_014_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                          //          .endofpacket
	);

	niosII_system_id_router_003 id_router_015 (
		.sink_ready         (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (solenoid_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                            //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset),                                      // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                    //       src.ready
		.src_valid          (id_router_015_src_valid),                                                    //          .valid
		.src_data           (id_router_015_src_data),                                                     //          .data
		.src_channel        (id_router_015_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                               //          .endofpacket
	);

	niosII_system_id_router_016 id_router_016 (
		.sink_ready         (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pwm_generator_0_avalon_slave_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                                 //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                                         //       src.ready
		.src_valid          (id_router_016_src_valid),                                                                         //          .valid
		.src_data           (id_router_016_src_data),                                                                          //          .data
		.src_channel        (id_router_016_src_channel),                                                                       //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                                 //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                                    //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (64),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.PKT_BURST_TYPE_H          (61),
		.PKT_BURST_TYPE_L          (60),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (54),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (86),
		.ST_CHANNEL_W              (17),
		.OUT_BYTE_CNT_H            (52),
		.OUT_BURSTWRAP_H           (56),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (altpll_0_c1_clk),                       //       cr0.clk
		.reset                 (nios2_0_jtag_debug_module_reset_reset), // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),               //     sink0.valid
		.sink0_data            (width_adapter_src_data),                //          .data
		.sink0_channel         (width_adapter_src_channel),             //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),       //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),         //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),               //          .ready
		.source0_valid         (burst_adapter_source0_valid),           //   source0.valid
		.source0_data          (burst_adapter_source0_data),            //          .data
		.source0_channel       (burst_adapter_source0_channel),         //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket),   //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),     //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)            //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (35),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (55),
		.PKT_BYTE_CNT_H            (44),
		.PKT_BYTE_CNT_L            (42),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (50),
		.PKT_BURST_SIZE_L          (48),
		.PKT_BURST_TYPE_H          (52),
		.PKT_BURST_TYPE_L          (51),
		.PKT_BURSTWRAP_H           (47),
		.PKT_BURSTWRAP_L           (45),
		.PKT_TRANS_COMPRESSED_READ (36),
		.PKT_TRANS_WRITE           (38),
		.PKT_TRANS_READ            (39),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (77),
		.ST_CHANNEL_W              (17),
		.OUT_BYTE_CNT_H            (42),
		.OUT_BURSTWRAP_H           (47),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter_001 (
		.clk                   (altpll_0_c1_clk),                         //       cr0.clk
		.reset                 (nios2_0_jtag_debug_module_reset_reset),   // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_n),                              // reset_in0.reset
		.reset_in1  (nios2_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (altpll_0_c1_clk),                       //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),        // reset_out.reset
		.reset_in2  (1'b0),                                  // (terminated)
		.reset_in3  (1'b0),                                  // (terminated)
		.reset_in4  (1'b0),                                  // (terminated)
		.reset_in5  (1'b0),                                  // (terminated)
		.reset_in6  (1'b0),                                  // (terminated)
		.reset_in7  (1'b0),                                  // (terminated)
		.reset_in8  (1'b0),                                  // (terminated)
		.reset_in9  (1'b0),                                  // (terminated)
		.reset_in10 (1'b0),                                  // (terminated)
		.reset_in11 (1'b0),                                  // (terminated)
		.reset_in12 (1'b0),                                  // (terminated)
		.reset_in13 (1'b0),                                  // (terminated)
		.reset_in14 (1'b0),                                  // (terminated)
		.reset_in15 (1'b0)                                   // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_n),                              // reset_in0.reset
		.reset_in1  (nios2_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_0),                                 //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),    // reset_out.reset
		.reset_in2  (1'b0),                                  // (terminated)
		.reset_in3  (1'b0),                                  // (terminated)
		.reset_in4  (1'b0),                                  // (terminated)
		.reset_in5  (1'b0),                                  // (terminated)
		.reset_in6  (1'b0),                                  // (terminated)
		.reset_in7  (1'b0),                                  // (terminated)
		.reset_in8  (1'b0),                                  // (terminated)
		.reset_in9  (1'b0),                                  // (terminated)
		.reset_in10 (1'b0),                                  // (terminated)
		.reset_in11 (1'b0),                                  // (terminated)
		.reset_in12 (1'b0),                                  // (terminated)
		.reset_in13 (1'b0),                                  // (terminated)
		.reset_in14 (1'b0),                                  // (terminated)
		.reset_in15 (1'b0)                                   // (terminated)
	);

	niosII_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (altpll_0_c1_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (altpll_0_c1_clk),                        //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (altpll_0_c1_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (clk_0),                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_006 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_007 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_008 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_009 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_010 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_011 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_012 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_013 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_014 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_015 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_003 rsp_xbar_demux_016 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (altpll_0_c1_clk),                       //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (crosser_001_out_ready),                 //     sink5.ready
		.sink5_valid          (crosser_001_out_valid),                 //          .valid
		.sink5_channel        (crosser_001_out_channel),               //          .channel
		.sink5_data           (crosser_001_out_data),                  //          .data
		.sink5_startofpacket  (crosser_001_out_startofpacket),         //          .startofpacket
		.sink5_endofpacket    (crosser_001_out_endofpacket),           //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (62),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (71),
		.IN_PKT_BYTE_CNT_L             (69),
		.IN_PKT_TRANS_COMPRESSED_READ  (63),
		.IN_PKT_BURSTWRAP_H            (74),
		.IN_PKT_BURSTWRAP_L            (72),
		.IN_PKT_BURST_SIZE_H           (77),
		.IN_PKT_BURST_SIZE_L           (75),
		.IN_PKT_RESPONSE_STATUS_H      (103),
		.IN_PKT_RESPONSE_STATUS_L      (102),
		.IN_PKT_TRANS_EXCLUSIVE        (68),
		.IN_PKT_BURST_TYPE_H           (79),
		.IN_PKT_BURST_TYPE_L           (78),
		.IN_ST_DATA_W                  (104),
		.OUT_PKT_ADDR_H                (44),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (53),
		.OUT_PKT_BYTE_CNT_L            (51),
		.OUT_PKT_TRANS_COMPRESSED_READ (45),
		.OUT_PKT_BURST_SIZE_H          (59),
		.OUT_PKT_BURST_SIZE_L          (57),
		.OUT_PKT_RESPONSE_STATUS_H     (85),
		.OUT_PKT_RESPONSE_STATUS_L     (84),
		.OUT_PKT_TRANS_EXCLUSIVE       (50),
		.OUT_PKT_BURST_TYPE_H          (61),
		.OUT_PKT_BURST_TYPE_L          (60),
		.OUT_ST_DATA_W                 (86),
		.ST_CHANNEL_W                  (17),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (altpll_0_c1_clk),                       //       clk.clk
		.reset                (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_mux_002_src_valid),            //      sink.valid
		.in_channel           (cmd_xbar_mux_002_src_channel),          //          .channel
		.in_startofpacket     (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.in_ready             (cmd_xbar_mux_002_src_ready),            //          .ready
		.in_data              (cmd_xbar_mux_002_src_data),             //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),         //       src.endofpacket
		.out_data             (width_adapter_src_data),                //          .data
		.out_channel          (width_adapter_src_channel),             //          .channel
		.out_valid            (width_adapter_src_valid),               //          .valid
		.out_ready            (width_adapter_src_ready),               //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),       //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (44),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (53),
		.IN_PKT_BYTE_CNT_L             (51),
		.IN_PKT_TRANS_COMPRESSED_READ  (45),
		.IN_PKT_BURSTWRAP_H            (56),
		.IN_PKT_BURSTWRAP_L            (54),
		.IN_PKT_BURST_SIZE_H           (59),
		.IN_PKT_BURST_SIZE_L           (57),
		.IN_PKT_RESPONSE_STATUS_H      (85),
		.IN_PKT_RESPONSE_STATUS_L      (84),
		.IN_PKT_TRANS_EXCLUSIVE        (50),
		.IN_PKT_BURST_TYPE_H           (61),
		.IN_PKT_BURST_TYPE_L           (60),
		.IN_ST_DATA_W                  (86),
		.OUT_PKT_ADDR_H                (62),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (71),
		.OUT_PKT_BYTE_CNT_L            (69),
		.OUT_PKT_TRANS_COMPRESSED_READ (63),
		.OUT_PKT_BURST_SIZE_H          (77),
		.OUT_PKT_BURST_SIZE_L          (75),
		.OUT_PKT_RESPONSE_STATUS_H     (103),
		.OUT_PKT_RESPONSE_STATUS_L     (102),
		.OUT_PKT_TRANS_EXCLUSIVE       (68),
		.OUT_PKT_BURST_TYPE_H          (79),
		.OUT_PKT_BURST_TYPE_L          (78),
		.OUT_ST_DATA_W                 (104),
		.ST_CHANNEL_W                  (17),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (altpll_0_c1_clk),                       //       clk.clk
		.reset                (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.in_valid             (id_router_002_src_valid),               //      sink.valid
		.in_channel           (id_router_002_src_channel),             //          .channel
		.in_startofpacket     (id_router_002_src_startofpacket),       //          .startofpacket
		.in_endofpacket       (id_router_002_src_endofpacket),         //          .endofpacket
		.in_ready             (id_router_002_src_ready),               //          .ready
		.in_data              (id_router_002_src_data),                //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_001_src_data),            //          .data
		.out_channel          (width_adapter_001_src_channel),         //          .channel
		.out_valid            (width_adapter_001_src_valid),           //          .valid
		.out_ready            (width_adapter_001_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (62),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (71),
		.IN_PKT_BYTE_CNT_L             (69),
		.IN_PKT_TRANS_COMPRESSED_READ  (63),
		.IN_PKT_BURSTWRAP_H            (74),
		.IN_PKT_BURSTWRAP_L            (72),
		.IN_PKT_BURST_SIZE_H           (77),
		.IN_PKT_BURST_SIZE_L           (75),
		.IN_PKT_RESPONSE_STATUS_H      (103),
		.IN_PKT_RESPONSE_STATUS_L      (102),
		.IN_PKT_TRANS_EXCLUSIVE        (68),
		.IN_PKT_BURST_TYPE_H           (79),
		.IN_PKT_BURST_TYPE_L           (78),
		.IN_ST_DATA_W                  (104),
		.OUT_PKT_ADDR_H                (35),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (44),
		.OUT_PKT_BYTE_CNT_L            (42),
		.OUT_PKT_TRANS_COMPRESSED_READ (36),
		.OUT_PKT_BURST_SIZE_H          (50),
		.OUT_PKT_BURST_SIZE_L          (48),
		.OUT_PKT_RESPONSE_STATUS_H     (76),
		.OUT_PKT_RESPONSE_STATUS_L     (75),
		.OUT_PKT_TRANS_EXCLUSIVE       (41),
		.OUT_PKT_BURST_TYPE_H          (52),
		.OUT_PKT_BURST_TYPE_L          (51),
		.OUT_ST_DATA_W                 (77),
		.ST_CHANNEL_W                  (17),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (altpll_0_c1_clk),                        //       clk.clk
		.reset                (nios2_0_jtag_debug_module_reset_reset),  // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src16_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src16_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src16_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src16_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_002_src_data),             //          .data
		.out_channel          (width_adapter_002_src_channel),          //          .channel
		.out_valid            (width_adapter_002_src_valid),            //          .valid
		.out_ready            (width_adapter_002_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (35),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (44),
		.IN_PKT_BYTE_CNT_L             (42),
		.IN_PKT_TRANS_COMPRESSED_READ  (36),
		.IN_PKT_BURSTWRAP_H            (47),
		.IN_PKT_BURSTWRAP_L            (45),
		.IN_PKT_BURST_SIZE_H           (50),
		.IN_PKT_BURST_SIZE_L           (48),
		.IN_PKT_RESPONSE_STATUS_H      (76),
		.IN_PKT_RESPONSE_STATUS_L      (75),
		.IN_PKT_TRANS_EXCLUSIVE        (41),
		.IN_PKT_BURST_TYPE_H           (52),
		.IN_PKT_BURST_TYPE_L           (51),
		.IN_ST_DATA_W                  (77),
		.OUT_PKT_ADDR_H                (62),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (71),
		.OUT_PKT_BYTE_CNT_L            (69),
		.OUT_PKT_TRANS_COMPRESSED_READ (63),
		.OUT_PKT_BURST_SIZE_H          (77),
		.OUT_PKT_BURST_SIZE_L          (75),
		.OUT_PKT_RESPONSE_STATUS_H     (103),
		.OUT_PKT_RESPONSE_STATUS_L     (102),
		.OUT_PKT_TRANS_EXCLUSIVE       (68),
		.OUT_PKT_BURST_TYPE_H          (79),
		.OUT_PKT_BURST_TYPE_L          (78),
		.OUT_ST_DATA_W                 (104),
		.ST_CHANNEL_W                  (17),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_003 (
		.clk                  (altpll_0_c1_clk),                       //       clk.clk
		.reset                (nios2_0_jtag_debug_module_reset_reset), // clk_reset.reset
		.in_valid             (id_router_016_src_valid),               //      sink.valid
		.in_channel           (id_router_016_src_channel),             //          .channel
		.in_startofpacket     (id_router_016_src_startofpacket),       //          .startofpacket
		.in_endofpacket       (id_router_016_src_endofpacket),         //          .endofpacket
		.in_ready             (id_router_016_src_ready),               //          .ready
		.in_data              (id_router_016_src_data),                //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_003_src_data),            //          .data
		.out_channel          (width_adapter_003_src_channel),         //          .channel
		.out_valid            (width_adapter_003_src_valid),           //          .valid
		.out_ready            (width_adapter_003_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (104),
		.BITS_PER_SYMBOL     (104),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (17),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (altpll_0_c1_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_0),                                 //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src5_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src5_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src5_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src5_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src5_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (104),
		.BITS_PER_SYMBOL     (104),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (17),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_0),                                 //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c1_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_005_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_005_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_005_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_005_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	niosII_system_irq_mapper irq_mapper (
		.clk           (altpll_0_c1_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_0_d_irq_irq)               //    sender.irq
	);

endmodule
